`ifndef CONSTANTS
`define CONSTANTS

// digital clock
    `define MODE_CLOCK 0
    `define MODE_TIMER 1
    `define MODE_ALARM 2

// edit time
    `define SELECT_NONE 0
    `define SELECT_SEC 1
    `define SELECT_MIN 2
    `define SELECT_HOUR 3

// 
    `define MEGA 1_000_000
    `define KILO 1_000
`endif
